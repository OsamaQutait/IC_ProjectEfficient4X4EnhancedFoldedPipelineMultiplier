*** SPICE deck for cell not{sch} from library Multiplier
*** Created on Fri Sep 01, 2023 18:51:13
*** Last revised on Fri Sep 08, 2023 10:21:34
*** Written on Fri Sep 08, 2023 10:21:39 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: not{sch}
Mnmos@0 out in gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd in out vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'not{sch}'
vdd vdd 0 DC 5V
v0 in 0 DC 5V pulse(0V 5V 0 0.1ns 0.1ns 10ns 20ns)
cload0 out 0 20fF
.tran 200ns
.include C:\Users\user\Downloads\C5_models.txt"
.END

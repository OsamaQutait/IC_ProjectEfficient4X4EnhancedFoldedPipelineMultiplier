*** SPICE deck for cell mux{sch} from library Multiplier
*** Created on Fri Sep 01, 2023 18:52:24
*** Last revised on Fri Sep 01, 2023 22:08:00
*** Written on Wed Sep 06, 2023 19:03:12 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Multiplier__not FROM CELL not{sch}
.SUBCKT Multiplier__not in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd in out vdd PMOS L=0.4U W=2U
.ENDS Multiplier__not

.global gnd vdd

*** TOP LEVEL CELL: mux{sch}
Mnmos@0 a sel out gnd NMOS L=0.4U W=2U
Mnmos@1 b net@29 out gnd NMOS L=0.4U W=2U
Mpmos@0 out net@29 a vdd PMOS L=0.4U W=2U
Mpmos@1 out sel b vdd PMOS L=0.4U W=2U
Xnot@0 sel net@29 Multiplier__not

* Spice Code nodes in cell cell 'mux{sch}'
vdd vdd 0 DC 5V
v1 a 0 DC 5V pulse(0V 5V 0 0.1ns 0.1ns 10ns 20ns)
v2 b 0 DC 5V pulse(0V 5V 0 0.1ns 0.1ns 10ns 40ns)
v3 sel 0 DC 5V pulse(0V 5V 0 0.1ns 0.1ns 10ns 80ns)
cload out 0 20fF
.tran 200ns
.include C:\Users\user\Downloads\C5_models.txt
.END

*** SPICE deck for cell xor{sch} from library Multiplier
*** Created on Fri Sep 01, 2023 18:52:10
*** Last revised on Fri Sep 08, 2023 10:08:29
*** Written on Fri Sep 08, 2023 10:08:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Multiplier__not FROM CELL not{sch}
.SUBCKT Multiplier__not in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.4U W=2U
Mpmos@0 vdd in out vdd PMOS L=0.4U W=2U
.ENDS Multiplier__not

.global gnd vdd

*** TOP LEVEL CELL: xor{sch}
Mnmos@0 a net@29 out gnd NMOS L=0.4U W=2U
Mnmos@1 net@16 b out gnd NMOS L=0.4U W=2U
Mpmos@0 out b a vdd PMOS L=0.4U W=2U
Mpmos@1 out net@29 net@16 vdd PMOS L=0.4U W=2U
Xnot@0 a net@16 Multiplier__not
Xnot@1 b net@29 Multiplier__not

* Spice Code nodes in cell cell 'xor{sch}'
vdd vdd 0 DC 5V
v0 a 0 DC 5V pulse(0V 5V 0 0.1ns 0.1ns 10ns 20ns)
v1 b 0 DC 5V pulse(0V 5V 0 0.1ns 0.1ns 10ns 40ns)
cload0 out 0 20fF
.tran 200ns
.include C:\Users\user\Downloads\C5_models.txt"
.END
